module top(
    input               i_clk,

    input       [4:0]   i_key,
    output      [3:0]   o_led,o_core_led,

    input               i_uart_rx,
    output              o_uart_tx,

    output              o_hdmi_clk_p,
    output              o_hdmi_clk_n,
    output      [2:0]   o_hdmi_d_p,
    output      [2:0]   o_hdmi_d_n,

    output      [13:0]  exter_io1
);
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			    测试时钟输入 	         /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
// 降低到hz，生成分频信号1hz A
logic [24:0] cnt;
always@(posedge i_clk)
    cnt <= cnt + 1;

logic clk_A ;
assign clk_A = cnt[24];

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 		        测试按键LED	            /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//现象：按键按下，对应的LED灭，否则 闪烁 

assign   o_led[0] = ~i_key[0] ? 1'd0 : cnt[23];
assign   o_led[1] = ~i_key[1] ? 1'd0 : cnt[23];
assign   o_led[2] = ~i_key[2] ? 1'd0 : cnt[23];
assign   o_led[3] = ~i_key[3] ? 1'd0 : cnt[23];

assign   o_core_led[0] = ~i_key[4]? 1'b0: cnt[23];
assign   o_core_led[1] = ~i_key[4]? 1'b0: cnt[23];
assign   o_core_led[2] = ~i_key[4]? 1'b0: cnt[23];
assign   o_core_led[3] = ~i_key[4]? 1'b0: cnt[23];


/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			    测试FLASH 	            /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//测试固化代码是否成功

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			    测试UART	            /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//回环测试
assign o_uart_tx = i_uart_rx;

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			    测试外部IO	            /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
assign exter_io1[0] = clk_A ;
assign exter_io1[1] = ~clk_A ;
assign exter_io1[2] = clk_A ;
assign exter_io1[3] = ~clk_A ;
assign exter_io1[4] = clk_A ;
assign exter_io1[5] = ~clk_A ;
assign exter_io1[6] = clk_A ;
assign exter_io1[7] = ~clk_A ;
assign exter_io1[8] = clk_A ;
assign exter_io1[9] = ~clk_A ;
assign exter_io1[10] = clk_A ;
assign exter_io1[11] = ~clk_A ;
assign exter_io1[12] = clk_A ;
assign exter_io1[13] = ~clk_A ;

/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
//////////////////// 			    测试HDMI	            /////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////

hdmi_colorbar_top hdmi_colorbar_top_m0(
	.sys_clk			(i_clk	 		),
	.sys_rst_n			(1'b1  			),
	.tmds_clk_p			(o_hdmi_clk_p	),
	.tmds_clk_n			(o_hdmi_clk_n	),
	.tmds_oen			(				),
	.tmds_data_p		(o_hdmi_d_p		),
	.tmds_data_n		(o_hdmi_d_n		)
);


endmodule 